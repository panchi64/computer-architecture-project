// Test Code
`timescale 1ns/1ns

module SOH_tb;

    reg [31:0] RB, PC;
    reg [11:0] imm12_I, imm12_S;
    reg [19:0] imm20;

    wire [31:0] N;

endmodule